class ahb_mtrxn extends uvm_sequence_item;
    // This file defines the AHB master transaction class
endclass: ahb_mtrxn